module cpu (
    
);

// Everything is in `cpu_datapath.sv`
    
endmodule