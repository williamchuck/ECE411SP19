module cpu_control (
    /// TODO: Consult Richard for the control interface.
);
    /// MARK: - Control word based on opcode (as outlined in the MP3 handout)
endmodule