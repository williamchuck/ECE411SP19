module hdu (
    /// TODO: Consult Richard for the HDU interface.
    output logic no_hazard
);

assign no_hazard = 1'd1;
    
endmodule