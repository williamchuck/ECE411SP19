module pc_register #(parameter width = 32)
(
    input clk,
    input load,
    input [width-1:0] in,
    output logic [width-1:0] out
);

logic [width-1:0] data;

/*
* PC needs to start at 0x60
 */
initial
begin
    data = 32'h00000060;
end

always_ff @(posedge clk)
begin
    if (load) begin
        data <= in;
    end
end

always_comb
begin
    out = data;
end

endmodule : pc_register
