module cpu (
    
);
    
endmodule