module fwu (
    /// TODO: Consult Richard for the FWU interface.
);
    
endmodule