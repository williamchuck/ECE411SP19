module hdu (
    /// TODO: Consult Richard for the HDU interface.
);
    
endmodule